//  Author  Lutz Filor
//  Date    04-13-2020
//  Email   lutz@pacbell.net
//  Phone   408-807-6915
//  ============================================================================
//
interface

